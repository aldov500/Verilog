library verilog;
use verilog.vl_types.all;
entity Example_03_05 is
end Example_03_05;
