library verilog;
use verilog.vl_types.all;
entity Example_04_03 is
end Example_04_03;
