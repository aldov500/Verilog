library verilog;
use verilog.vl_types.all;
entity Example_06_03 is
end Example_06_03;
