library verilog;
use verilog.vl_types.all;
entity Router is
end Router;
