library verilog;
use verilog.vl_types.all;
entity Example_03_07_02 is
end Example_03_07_02;
