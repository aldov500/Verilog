library verilog;
use verilog.vl_types.all;
entity Example_04_04 is
end Example_04_04;
