library verilog;
use verilog.vl_types.all;
entity example33 is
end example33;
