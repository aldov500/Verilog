library verilog;
use verilog.vl_types.all;
entity PkgB is
end PkgB;
