library verilog;
use verilog.vl_types.all;
entity Example_02_03 is
end Example_02_03;
