library verilog;
use verilog.vl_types.all;
entity Example_05_02 is
end Example_05_02;
