library verilog;
use verilog.vl_types.all;
entity Example_02_02 is
end Example_02_02;
