library verilog;
use verilog.vl_types.all;
entity Example_04_01 is
end Example_04_01;
