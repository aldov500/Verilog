library verilog;
use verilog.vl_types.all;
entity EnvPkg is
end EnvPkg;
