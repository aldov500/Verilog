library verilog;
use verilog.vl_types.all;
entity TaskPkg is
end TaskPkg;
