library verilog;
use verilog.vl_types.all;
entity example31 is
end example31;
