library verilog;
use verilog.vl_types.all;
entity Example_03_07_04 is
end Example_03_07_04;
