library verilog;
use verilog.vl_types.all;
entity Example_06_06 is
end Example_06_06;
