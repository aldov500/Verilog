library verilog;
use verilog.vl_types.all;
entity Example_03_07_03 is
end Example_03_07_03;
