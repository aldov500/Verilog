library verilog;
use verilog.vl_types.all;
entity example30 is
end example30;
