library verilog;
use verilog.vl_types.all;
entity Example_03_03 is
end Example_03_03;
