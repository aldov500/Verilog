library verilog;
use verilog.vl_types.all;
entity Example_05_04_02 is
end Example_05_04_02;
