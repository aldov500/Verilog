library verilog;
use verilog.vl_types.all;
entity Example_03_06_01 is
end Example_03_06_01;
