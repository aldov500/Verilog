library verilog;
use verilog.vl_types.all;
entity PkgA is
end PkgA;
