library verilog;
use verilog.vl_types.all;
entity Example_03_01 is
end Example_03_01;
